module pkkg;
function [3:0] addd;
input [3:0] a,b;
begin
  addd = a+b;
end
endfunction
endmodule
